// module of NEOcalculator
timeunit 1ns; timeprecision 10ps;

module NEOcalculator #(
    parameter N = 16,  // N-bits wide
    parameter M = 32  // M locations
    )(
    input logic Clk,
    input logic reset,
    input logic signed [N-1:0] rdata,
    output logic [$clog2(M)-1:0] raddr,
    output logic [$clog2(M)-1:0] waddr,
    output logic signed [N-1:0] wdata,
    output logic ready
);



logic signed [N-1:0] xn_prev, xn_curr;
logic [$clog2(M):0] counter;

always_ff @(posedge Clk, negedge reset) begin
    if (!reset) begin
        counter <= '0;
        xn_prev <= '0;
        xn_curr <= '0;
        ready <= '0;

    end else begin
        // Simple processing: shift data through registers
    xn_curr <= rdata;
    xn_prev <= xn_curr;   


    if (counter >= (M + 2)) begin
        counter <= counter;     // hold
        ready   <= 1'b0;

    
    end else if (counter == (M + 1)) begin
        counter <= counter + 1;
        ready   <= 1'b1;


    end else begin
        counter <= counter + 1;
    end

    end
end

always_comb begin
    if (counter >= 2) begin
        waddr = counter - 2;
    end else begin
        waddr = '0;
    end
    
    if (counter >= M-1) begin
    raddr = M-1;
    end else begin
    raddr = counter;
    end

    wdata = xn_curr * xn_curr - rdata * xn_prev;
end

endmodule