// module of Toplevel
